/*
* Copyright (c) 2024 Your Name
* SPDX-License-Identifier: Apache-2.0
*/
`default_nettype none
 
module EjemploSUMADOR1BIT (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
 wire s1, c1, s2;
  // instance
  C_XOR U1(.OUT(s1),    .A(ui_in[0]),  .B(ui_in[1])); // es la compuerta 1 
  C_AND U2(.OUT(c1),    .A(ui_in[0]),  .B(ui_in[1])); // la sintaxis es salida entrada entrada
  C_XOR U3(.OUT(uo_out[0]),  .A(s1), .B(ui_in[2]));
  C_AND U4(.OUT(s2),    .A(s1), .B(ui_in[2]));
  C_XOR U5(.OUT(uo_out[1]), .A(s2), .B(c1));
  
  // All output pins must be assigned. If not used, assign to 0.
  assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;
 
  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};
endmodule
